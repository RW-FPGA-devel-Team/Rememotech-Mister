    r(0) := x"f3";
    r(1) := x"31";
    r(2) := x"00";
    r(3) := x"ff";
    r(4) := x"cd";
    r(5) := x"45";
    r(6) := x"00";
    r(7) := x"db";
    r(8) := x"c5";
    r(9) := x"f5";
    r(10) := x"cb";
    r(11) := x"57";
    r(12) := x"cc";
    r(13) := x"8a";
    r(14) := x"00";
    r(15) := x"f1";
    r(16) := x"f5";
    r(17) := x"cb";
    r(18) := x"4f";
    r(19) := x"cc";
    r(20) := x"36";
    r(21) := x"01";
    r(22) := x"f1";
    r(23) := x"cb";
    r(24) := x"47";
    r(25) := x"cc";
    r(26) := x"40";
    r(27) := x"01";
    r(28) := x"3e";
    r(29) := x"08";
    r(30) := x"d3";
    r(31) := x"d0";
    r(32) := x"21";
    r(33) := x"00";
    r(34) := x"60";
    r(35) := x"11";
    r(36) := x"3d";
    r(37) := x"00";
    r(38) := x"06";
    r(39) := x"08";
    r(40) := x"1a";
    r(41) := x"be";
    r(42) := x"20";
    r(43) := x"0c";
    r(44) := x"13";
    r(45) := x"23";
    r(46) := x"10";
    r(47) := x"f8";
    r(48) := x"af";
    r(49) := x"d3";
    r(50) := x"c0";
    r(51) := x"d3";
    r(52) := x"c1";
    r(53) := x"c3";
    r(54) := x"08";
    r(55) := x"60";
    r(56) := x"3e";
    r(57) := x"ff";
    r(58) := x"c3";
    r(59) := x"5d";
    r(60) := x"02";
    r(61) := x"52";
    r(62) := x"45";
    r(63) := x"4d";
    r(64) := x"4f";
    r(65) := x"4e";
    r(66) := x"35";
    r(67) := x"31";
    r(68) := x"32";
    r(69) := x"3e";
    r(70) := x"0c";
    r(71) := x"d3";
    r(72) := x"38";
    r(73) := x"af";
    r(74) := x"d3";
    r(75) := x"39";
    r(76) := x"3e";
    r(77) := x"0d";
    r(78) := x"d3";
    r(79) := x"38";
    r(80) := x"af";
    r(81) := x"d3";
    r(82) := x"39";
    r(83) := x"3e";
    r(84) := x"0e";
    r(85) := x"d3";
    r(86) := x"38";
    r(87) := x"af";
    r(88) := x"d3";
    r(89) := x"39";
    r(90) := x"3e";
    r(91) := x"0f";
    r(92) := x"d3";
    r(93) := x"38";
    r(94) := x"af";
    r(95) := x"d3";
    r(96) := x"39";
    r(97) := x"3e";
    r(98) := x"0a";
    r(99) := x"d3";
    r(100) := x"38";
    r(101) := x"af";
    r(102) := x"d3";
    r(103) := x"39";
    r(104) := x"3e";
    r(105) := x"1f";
    r(106) := x"d3";
    r(107) := x"38";
    r(108) := x"af";
    r(109) := x"d3";
    r(110) := x"39";
    r(111) := x"3e";
    r(112) := x"20";
    r(113) := x"d3";
    r(114) := x"32";
    r(115) := x"3e";
    r(116) := x"07";
    r(117) := x"d3";
    r(118) := x"33";
    r(119) := x"21";
    r(120) := x"00";
    r(121) := x"e0";
    r(122) := x"01";
    r(123) := x"00";
    r(124) := x"10";
    r(125) := x"7c";
    r(126) := x"d3";
    r(127) := x"31";
    r(128) := x"7d";
    r(129) := x"d3";
    r(130) := x"30";
    r(131) := x"23";
    r(132) := x"0b";
    r(133) := x"78";
    r(134) := x"b1";
    r(135) := x"20";
    r(136) := x"f4";
    r(137) := x"c9";
    r(138) := x"3e";
    r(139) := x"20";
    r(140) := x"d3";
    r(141) := x"c1";
    r(142) := x"cd";
    r(143) := x"5e";
    r(144) := x"01";
    r(145) := x"3e";
    r(146) := x"0a";
    r(147) := x"cd";
    r(148) := x"ac";
    r(149) := x"01";
    r(150) := x"3e";
    r(151) := x"09";
    r(152) := x"cd";
    r(153) := x"ac";
    r(154) := x"01";
    r(155) := x"21";
    r(156) := x"80";
    r(157) := x"00";
    r(158) := x"22";
    r(159) := x"20";
    r(160) := x"fe";
    r(161) := x"21";
    r(162) := x"00";
    r(163) := x"00";
    r(164) := x"22";
    r(165) := x"22";
    r(166) := x"fe";
    r(167) := x"3e";
    r(168) := x"01";
    r(169) := x"06";
    r(170) := x"07";
    r(171) := x"c5";
    r(172) := x"f5";
    r(173) := x"cb";
    r(174) := x"27";
    r(175) := x"cb";
    r(176) := x"27";
    r(177) := x"d3";
    r(178) := x"d1";
    r(179) := x"3e";
    r(180) := x"f0";
    r(181) := x"32";
    r(182) := x"aa";
    r(183) := x"8a";
    r(184) := x"3e";
    r(185) := x"aa";
    r(186) := x"32";
    r(187) := x"aa";
    r(188) := x"8a";
    r(189) := x"3e";
    r(190) := x"55";
    r(191) := x"32";
    r(192) := x"55";
    r(193) := x"85";
    r(194) := x"3e";
    r(195) := x"80";
    r(196) := x"32";
    r(197) := x"aa";
    r(198) := x"8a";
    r(199) := x"3e";
    r(200) := x"aa";
    r(201) := x"32";
    r(202) := x"aa";
    r(203) := x"8a";
    r(204) := x"3e";
    r(205) := x"55";
    r(206) := x"32";
    r(207) := x"55";
    r(208) := x"85";
    r(209) := x"3e";
    r(210) := x"30";
    r(211) := x"32";
    r(212) := x"00";
    r(213) := x"80";
    r(214) := x"06";
    r(215) := x"ff";
    r(216) := x"10";
    r(217) := x"fe";
    r(218) := x"3a";
    r(219) := x"00";
    r(220) := x"80";
    r(221) := x"cb";
    r(222) := x"7f";
    r(223) := x"28";
    r(224) := x"f9";
    r(225) := x"f1";
    r(226) := x"f5";
    r(227) := x"06";
    r(228) := x"04";
    r(229) := x"4f";
    r(230) := x"cb";
    r(231) := x"21";
    r(232) := x"cb";
    r(233) := x"21";
    r(234) := x"c5";
    r(235) := x"11";
    r(236) := x"00";
    r(237) := x"80";
    r(238) := x"79";
    r(239) := x"d3";
    r(240) := x"c0";
    r(241) := x"d3";
    r(242) := x"d1";
    r(243) := x"06";
    r(244) := x"20";
    r(245) := x"c5";
    r(246) := x"21";
    r(247) := x"00";
    r(248) := x"fc";
    r(249) := x"cd";
    r(250) := x"e2";
    r(251) := x"01";
    r(252) := x"01";
    r(253) := x"00";
    r(254) := x"02";
    r(255) := x"21";
    r(256) := x"00";
    r(257) := x"fc";
    r(258) := x"3e";
    r(259) := x"aa";
    r(260) := x"32";
    r(261) := x"aa";
    r(262) := x"8a";
    r(263) := x"3e";
    r(264) := x"55";
    r(265) := x"32";
    r(266) := x"55";
    r(267) := x"85";
    r(268) := x"3e";
    r(269) := x"a0";
    r(270) := x"32";
    r(271) := x"aa";
    r(272) := x"8a";
    r(273) := x"7e";
    r(274) := x"12";
    r(275) := x"1a";
    r(276) := x"be";
    r(277) := x"20";
    r(278) := x"fc";
    r(279) := x"23";
    r(280) := x"13";
    r(281) := x"0b";
    r(282) := x"78";
    r(283) := x"b1";
    r(284) := x"20";
    r(285) := x"e4";
    r(286) := x"2a";
    r(287) := x"20";
    r(288) := x"fe";
    r(289) := x"23";
    r(290) := x"22";
    r(291) := x"20";
    r(292) := x"fe";
    r(293) := x"c1";
    r(294) := x"10";
    r(295) := x"cd";
    r(296) := x"c1";
    r(297) := x"0c";
    r(298) := x"10";
    r(299) := x"be";
    r(300) := x"f1";
    r(301) := x"3c";
    r(302) := x"c1";
    r(303) := x"05";
    r(304) := x"c2";
    r(305) := x"ab";
    r(306) := x"00";
    r(307) := x"c3";
    r(308) := x"a8";
    r(309) := x"01";
    r(310) := x"3e";
    r(311) := x"10";
    r(312) := x"d3";
    r(313) := x"c1";
    r(314) := x"06";
    r(315) := x"08";
    r(316) := x"3e";
    r(317) := x"04";
    r(318) := x"18";
    r(319) := x"07";
    r(320) := x"af";
    r(321) := x"d3";
    r(322) := x"c1";
    r(323) := x"06";
    r(324) := x"14";
    r(325) := x"3e";
    r(326) := x"0c";
    r(327) := x"c5";
    r(328) := x"d3";
    r(329) := x"c0";
    r(330) := x"d3";
    r(331) := x"d1";
    r(332) := x"d3";
    r(333) := x"d0";
    r(334) := x"21";
    r(335) := x"00";
    r(336) := x"80";
    r(337) := x"11";
    r(338) := x"00";
    r(339) := x"40";
    r(340) := x"01";
    r(341) := x"00";
    r(342) := x"40";
    r(343) := x"ed";
    r(344) := x"b0";
    r(345) := x"c1";
    r(346) := x"3c";
    r(347) := x"10";
    r(348) := x"ea";
    r(349) := x"c9";
    r(350) := x"3e";
    r(351) := x"3e";
    r(352) := x"d3";
    r(353) := x"d4";
    r(354) := x"06";
    r(355) := x"0a";
    r(356) := x"3e";
    r(357) := x"ff";
    r(358) := x"d3";
    r(359) := x"d6";
    r(360) := x"db";
    r(361) := x"d4";
    r(362) := x"cb";
    r(363) := x"7f";
    r(364) := x"28";
    r(365) := x"fa";
    r(366) := x"10";
    r(367) := x"f4";
    r(368) := x"3e";
    r(369) := x"be";
    r(370) := x"d3";
    r(371) := x"d4";
    r(372) := x"06";
    r(373) := x"ff";
    r(374) := x"c5";
    r(375) := x"af";
    r(376) := x"cd";
    r(377) := x"1d";
    r(378) := x"02";
    r(379) := x"c1";
    r(380) := x"fe";
    r(381) := x"01";
    r(382) := x"28";
    r(383) := x"07";
    r(384) := x"10";
    r(385) := x"f4";
    r(386) := x"3e";
    r(387) := x"01";
    r(388) := x"c3";
    r(389) := x"5d";
    r(390) := x"02";
    r(391) := x"01";
    r(392) := x"e8";
    r(393) := x"03";
    r(394) := x"c5";
    r(395) := x"3e";
    r(396) := x"37";
    r(397) := x"cd";
    r(398) := x"1d";
    r(399) := x"02";
    r(400) := x"3e";
    r(401) := x"29";
    r(402) := x"cd";
    r(403) := x"1d";
    r(404) := x"02";
    r(405) := x"c1";
    r(406) := x"a7";
    r(407) := x"28";
    r(408) := x"0a";
    r(409) := x"0b";
    r(410) := x"78";
    r(411) := x"b1";
    r(412) := x"20";
    r(413) := x"ec";
    r(414) := x"3e";
    r(415) := x"02";
    r(416) := x"c3";
    r(417) := x"5d";
    r(418) := x"02";
    r(419) := x"3e";
    r(420) := x"80";
    r(421) := x"d3";
    r(422) := x"d4";
    r(423) := x"c9";
    r(424) := x"af";
    r(425) := x"d3";
    r(426) := x"d4";
    r(427) := x"c9";
    r(428) := x"06";
    r(429) := x"0a";
    r(430) := x"c5";
    r(431) := x"cd";
    r(432) := x"1d";
    r(433) := x"02";
    r(434) := x"c1";
    r(435) := x"a7";
    r(436) := x"28";
    r(437) := x"08";
    r(438) := x"05";
    r(439) := x"28";
    r(440) := x"26";
    r(441) := x"cd";
    r(442) := x"50";
    r(443) := x"02";
    r(444) := x"18";
    r(445) := x"f0";
    r(446) := x"06";
    r(447) := x"0a";
    r(448) := x"cd";
    r(449) := x"50";
    r(450) := x"02";
    r(451) := x"fe";
    r(452) := x"fe";
    r(453) := x"28";
    r(454) := x"04";
    r(455) := x"10";
    r(456) := x"f5";
    r(457) := x"18";
    r(458) := x"14";
    r(459) := x"06";
    r(460) := x"10";
    r(461) := x"21";
    r(462) := x"00";
    r(463) := x"fe";
    r(464) := x"cd";
    r(465) := x"50";
    r(466) := x"02";
    r(467) := x"77";
    r(468) := x"23";
    r(469) := x"10";
    r(470) := x"f9";
    r(471) := x"cd";
    r(472) := x"50";
    r(473) := x"02";
    r(474) := x"cd";
    r(475) := x"50";
    r(476) := x"02";
    r(477) := x"af";
    r(478) := x"c9";
    r(479) := x"3e";
    r(480) := x"ff";
    r(481) := x"c9";
    r(482) := x"d5";
    r(483) := x"e5";
    r(484) := x"ed";
    r(485) := x"5b";
    r(486) := x"20";
    r(487) := x"fe";
    r(488) := x"2a";
    r(489) := x"22";
    r(490) := x"fe";
    r(491) := x"65";
    r(492) := x"6a";
    r(493) := x"53";
    r(494) := x"1e";
    r(495) := x"00";
    r(496) := x"cb";
    r(497) := x"22";
    r(498) := x"cb";
    r(499) := x"15";
    r(500) := x"cb";
    r(501) := x"14";
    r(502) := x"3e";
    r(503) := x"11";
    r(504) := x"cd";
    r(505) := x"23";
    r(506) := x"02";
    r(507) := x"06";
    r(508) := x"ff";
    r(509) := x"cd";
    r(510) := x"50";
    r(511) := x"02";
    r(512) := x"fe";
    r(513) := x"fe";
    r(514) := x"28";
    r(515) := x"07";
    r(516) := x"10";
    r(517) := x"f7";
    r(518) := x"3e";
    r(519) := x"03";
    r(520) := x"c3";
    r(521) := x"5d";
    r(522) := x"02";
    r(523) := x"01";
    r(524) := x"d7";
    r(525) := x"00";
    r(526) := x"e1";
    r(527) := x"e5";
    r(528) := x"ed";
    r(529) := x"78";
    r(530) := x"ed";
    r(531) := x"b2";
    r(532) := x"ed";
    r(533) := x"b2";
    r(534) := x"ed";
    r(535) := x"78";
    r(536) := x"db";
    r(537) := x"d6";
    r(538) := x"e1";
    r(539) := x"d1";
    r(540) := x"c9";
    r(541) := x"21";
    r(542) := x"00";
    r(543) := x"00";
    r(544) := x"11";
    r(545) := x"00";
    r(546) := x"00";
    r(547) := x"f5";
    r(548) := x"cd";
    r(549) := x"50";
    r(550) := x"02";
    r(551) := x"f1";
    r(552) := x"f6";
    r(553) := x"40";
    r(554) := x"cd";
    r(555) := x"52";
    r(556) := x"02";
    r(557) := x"7c";
    r(558) := x"cd";
    r(559) := x"52";
    r(560) := x"02";
    r(561) := x"7d";
    r(562) := x"cd";
    r(563) := x"52";
    r(564) := x"02";
    r(565) := x"7a";
    r(566) := x"cd";
    r(567) := x"52";
    r(568) := x"02";
    r(569) := x"7b";
    r(570) := x"cd";
    r(571) := x"52";
    r(572) := x"02";
    r(573) := x"3e";
    r(574) := x"95";
    r(575) := x"cd";
    r(576) := x"52";
    r(577) := x"02";
    r(578) := x"cd";
    r(579) := x"50";
    r(580) := x"02";
    r(581) := x"06";
    r(582) := x"0a";
    r(583) := x"cd";
    r(584) := x"50";
    r(585) := x"02";
    r(586) := x"cb";
    r(587) := x"7f";
    r(588) := x"c8";
    r(589) := x"10";
    r(590) := x"f8";
    r(591) := x"c9";
    r(592) := x"3e";
    r(593) := x"ff";
    r(594) := x"d3";
    r(595) := x"d6";
    r(596) := x"db";
    r(597) := x"d4";
    r(598) := x"cb";
    r(599) := x"7f";
    r(600) := x"28";
    r(601) := x"fa";
    r(602) := x"db";
    r(603) := x"d6";
    r(604) := x"c9";
    r(605) := x"d3";
    r(606) := x"c0";
    r(607) := x"3e";
    r(608) := x"ee";
    r(609) := x"d3";
    r(610) := x"c1";
    r(611) := x"18";
    r(612) := x"fe";
    r(613) := x"5b";
    r(614) := x"20";
    r(615) := x"fe";
    r(616) := x"2a";
    r(617) := x"22";
    r(618) := x"fe";
    r(619) := x"65";
    r(620) := x"6a";
    r(621) := x"53";
    r(622) := x"1e";
    r(623) := x"00";
    r(624) := x"cb";
    r(625) := x"22";
    r(626) := x"cb";
    r(627) := x"15";
    r(628) := x"cb";
    r(629) := x"14";
    r(630) := x"3e";
    r(631) := x"11";
    r(632) := x"cd";
    r(633) := x"23";
    r(634) := x"02";
    r(635) := x"06";
    r(636) := x"ff";
    r(637) := x"cd";
    r(638) := x"50";
    r(639) := x"02";
