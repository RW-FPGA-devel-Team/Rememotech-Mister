--
-- mon_prom_alpha.vhd - Alpha character generator
--
-- This is the 80 column character set.
-- The first row of each of the 256 characters is stored,
-- then the next row of each, etc..
-- In this way, addressing is row&char (no multiply by 10 needed)
--
-- This is a synchronous implementation
--

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity mon_prom_alpha is
  port
    (
    clk  : in  std_logic;
    addr : in  std_logic_vector(11 downto 0);
    q    : out std_logic_vector(07 downto 0)
    );
end mon_prom_alpha;

architecture behavior of mon_prom_alpha is

  type rom_type is array (0 to 2559) of std_logic_vector(7 downto 0);

  function init_rom return rom_type is
    variable r : rom_type := (others => (others => 'X'));
  begin
    r(   0) := "00000000";
    r(   1) := "00000000";
    r(   2) := "00000000";
    r(   3) := "00000000";
    r(   4) := "00000000";
    r(   5) := "00000000";
    r(   6) := "00000000";
    r(   7) := "00000000";
    r(   8) := "00000000";
    r(   9) := "00000000";
    r(  10) := "00000000";
    r(  11) := "00000000";
    r(  12) := "00000000";
    r(  13) := "00000000";
    r(  14) := "00000000";
    r(  15) := "00000000";
    r(  16) := "00000000";
    r(  17) := "00000000";
    r(  18) := "00000000";
    r(  19) := "00000000";
    r(  20) := "00000000";
    r(  21) := "00000000";
    r(  22) := "00000000";
    r(  23) := "00000000";
    r(  24) := "00000000";
    r(  25) := "00000000";
    r(  26) := "00000000";
    r(  27) := "00000000";
    r(  28) := "00000000";
    r(  29) := "00000000";
    r(  30) := "00000000";
    r(  31) := "00000000";
    r(  32) := "00000000";
    r(  33) := "00000000";
    r(  34) := "00000000";
    r(  35) := "00000000";
    r(  36) := "00000000";
    r(  37) := "00000000";
    r(  38) := "00000000";
    r(  39) := "00000000";
    r(  40) := "00000000";
    r(  41) := "00000000";
    r(  42) := "00000000";
    r(  43) := "00000000";
    r(  44) := "00000000";
    r(  45) := "00000000";
    r(  46) := "00000000";
    r(  47) := "00000000";
    r(  48) := "00000000";
    r(  49) := "00000000";
    r(  50) := "00000000";
    r(  51) := "00000000";
    r(  52) := "00000000";
    r(  53) := "00000000";
    r(  54) := "00000000";
    r(  55) := "00000000";
    r(  56) := "00000000";
    r(  57) := "00000000";
    r(  58) := "00000000";
    r(  59) := "00000000";
    r(  60) := "00000000";
    r(  61) := "00000000";
    r(  62) := "00000000";
    r(  63) := "00000000";
    r(  64) := "00000000";
    r(  65) := "00000000";
    r(  66) := "00000000";
    r(  67) := "00000000";
    r(  68) := "00000000";
    r(  69) := "00000000";
    r(  70) := "00000000";
    r(  71) := "00000000";
    r(  72) := "00000000";
    r(  73) := "00000000";
    r(  74) := "00000000";
    r(  75) := "00000000";
    r(  76) := "00000000";
    r(  77) := "00000000";
    r(  78) := "00000000";
    r(  79) := "00000000";
    r(  80) := "00000000";
    r(  81) := "00000000";
    r(  82) := "00000000";
    r(  83) := "00000000";
    r(  84) := "00000000";
    r(  85) := "00000000";
    r(  86) := "00000000";
    r(  87) := "00000000";
    r(  88) := "00000000";
    r(  89) := "00000000";
    r(  90) := "00000000";
    r(  91) := "00000000";
    r(  92) := "00000000";
    r(  93) := "00000000";
    r(  94) := "00000000";
    r(  95) := "00000000";
    r(  96) := "00000000";
    r(  97) := "00000000";
    r(  98) := "00000000";
    r(  99) := "00000000";
    r( 100) := "00000000";
    r( 101) := "00000000";
    r( 102) := "00000000";
    r( 103) := "00000000";
    r( 104) := "00000000";
    r( 105) := "00000000";
    r( 106) := "00000000";
    r( 107) := "00000000";
    r( 108) := "00000000";
    r( 109) := "00000000";
    r( 110) := "00000000";
    r( 111) := "00000000";
    r( 112) := "00000000";
    r( 113) := "00000000";
    r( 114) := "00000000";
    r( 115) := "00000000";
    r( 116) := "00000000";
    r( 117) := "00000000";
    r( 118) := "00000000";
    r( 119) := "00000000";
    r( 120) := "00000000";
    r( 121) := "00000000";
    r( 122) := "00000000";
    r( 123) := "00000000";
    r( 124) := "00000000";
    r( 125) := "00000000";
    r( 126) := "00000000";
    r( 127) := "00000000";
    r( 128) := "00000000";
    r( 129) := "00011000";
    r( 130) := "00011000";
    r( 131) := "00011000";
    r( 132) := "00000000";
    r( 133) := "00000000";
    r( 134) := "00011000";
    r( 135) := "00011000";
    r( 136) := "00011000";
    r( 137) := "00000000";
    r( 138) := "00011000";
    r( 139) := "00000000";
    r( 140) := "00000000";
    r( 141) := "00000000";
    r( 142) := "00000000";
    r( 143) := "00000000";
    r( 144) := "00100100";
    r( 145) := "00000000";
    r( 146) := "00000000";
    r( 147) := "00000000";
    r( 148) := "00000000";
    r( 149) := "00000000";
    r( 150) := "00100100";
    r( 151) := "00000000";
    r( 152) := "00000000";
    r( 153) := "00000000";
    r( 154) := "00000000";
    r( 155) := "00000000";
    r( 156) := "00000000";
    r( 157) := "00000000";
    r( 158) := "00000000";
    r( 159) := "00111100";
    r( 160) := "00000000";
    r( 161) := "00000000";
    r( 162) := "00000000";
    r( 163) := "00000000";
    r( 164) := "00000000";
    r( 165) := "00000000";
    r( 166) := "00000000";
    r( 167) := "00000000";
    r( 168) := "00000000";
    r( 169) := "00000000";
    r( 170) := "00000000";
    r( 171) := "00000000";
    r( 172) := "00000000";
    r( 173) := "00000000";
    r( 174) := "00000000";
    r( 175) := "00000000";
    r( 176) := "00000000";
    r( 177) := "00000000";
    r( 178) := "00000000";
    r( 179) := "00000000";
    r( 180) := "00000000";
    r( 181) := "00000000";
    r( 182) := "00000000";
    r( 183) := "00000000";
    r( 184) := "00000000";
    r( 185) := "00000000";
    r( 186) := "00000000";
    r( 187) := "00000000";
    r( 188) := "00000000";
    r( 189) := "00000000";
    r( 190) := "00000000";
    r( 191) := "00000000";
    r( 192) := "00000000";
    r( 193) := "00000000";
    r( 194) := "00000000";
    r( 195) := "00000000";
    r( 196) := "00000000";
    r( 197) := "00000000";
    r( 198) := "00000000";
    r( 199) := "00000000";
    r( 200) := "00000000";
    r( 201) := "00000000";
    r( 202) := "00000000";
    r( 203) := "00000000";
    r( 204) := "00000000";
    r( 205) := "00000000";
    r( 206) := "00000000";
    r( 207) := "00000000";
    r( 208) := "00000000";
    r( 209) := "00000000";
    r( 210) := "00000000";
    r( 211) := "00000000";
    r( 212) := "00000000";
    r( 213) := "00000000";
    r( 214) := "00000000";
    r( 215) := "00000000";
    r( 216) := "00000000";
    r( 217) := "00000000";
    r( 218) := "00000000";
    r( 219) := "00000000";
    r( 220) := "00000000";
    r( 221) := "00000000";
    r( 222) := "00000000";
    r( 223) := "00000000";
    r( 224) := "00000000";
    r( 225) := "00000000";
    r( 226) := "00000000";
    r( 227) := "00000000";
    r( 228) := "00000000";
    r( 229) := "00000000";
    r( 230) := "00000000";
    r( 231) := "00000000";
    r( 232) := "00000000";
    r( 233) := "00000000";
    r( 234) := "00000000";
    r( 235) := "00000000";
    r( 236) := "00000000";
    r( 237) := "00000000";
    r( 238) := "00000000";
    r( 239) := "00000000";
    r( 240) := "00000000";
    r( 241) := "00000000";
    r( 242) := "00000000";
    r( 243) := "00000000";
    r( 244) := "00000000";
    r( 245) := "00000000";
    r( 246) := "00000000";
    r( 247) := "00000000";
    r( 248) := "00000000";
    r( 249) := "00000000";
    r( 250) := "00000000";
    r( 251) := "00000000";
    r( 252) := "00000000";
    r( 253) := "00000000";
    r( 254) := "00000000";
    r( 255) := "00000000";
    r( 256) := "00000000";
    r( 257) := "00000000";
    r( 258) := "00011000";
    r( 259) := "00111100";
    r( 260) := "11111110";
    r( 261) := "11111110";
    r( 262) := "00000100";
    r( 263) := "00010000";
    r( 264) := "00001000";
    r( 265) := "00010000";
    r( 266) := "00010000";
    r( 267) := "00010000";
    r( 268) := "10010010";
    r( 269) := "00000010";
    r( 270) := "00000010";
    r( 271) := "00000000";
    r( 272) := "01101100";
    r( 273) := "00010000";
    r( 274) := "00010000";
    r( 275) := "00010000";
    r( 276) := "01111100";
    r( 277) := "00000000";
    r( 278) := "00100000";
    r( 279) := "00000000";
    r( 280) := "00011000";
    r( 281) := "00001000";
    r( 282) := "00010000";
    r( 283) := "00010000";
    r( 284) := "00000000";
    r( 285) := "00000000";
    r( 286) := "00000000";
    r( 287) := "00000000";
    r( 288) := "00000000";
    r( 289) := "00001000";
    r( 290) := "00100100";
    r( 291) := "00100100";
    r( 292) := "00001000";
    r( 293) := "00000000";
    r( 294) := "00110000";
    r( 295) := "00000100";
    r( 296) := "00000100";
    r( 297) := "00100000";
    r( 298) := "00001000";
    r( 299) := "00000000";
    r( 300) := "00000000";
    r( 301) := "00000000";
    r( 302) := "00000000";
    r( 303) := "00000000";
    r( 304) := "00111100";
    r( 305) := "00001000";
    r( 306) := "00111100";
    r( 307) := "00111100";
    r( 308) := "00000100";
    r( 309) := "01111100";
    r( 310) := "00011100";
    r( 311) := "01111110";
    r( 312) := "00111100";
    r( 313) := "00111100";
    r( 314) := "00000000";
    r( 315) := "00000000";
    r( 316) := "00000100";
    r( 317) := "00000000";
    r( 318) := "00100000";
    r( 319) := "00111100";
    r( 320) := "00011100";
    r( 321) := "00011000";
    r( 322) := "01111100";
    r( 323) := "00111100";
    r( 324) := "01111100";
    r( 325) := "01111110";
    r( 326) := "01111110";
    r( 327) := "00111100";
    r( 328) := "01000010";
    r( 329) := "00011100";
    r( 330) := "00001110";
    r( 331) := "01000010";
    r( 332) := "01000000";
    r( 333) := "01000010";
    r( 334) := "01000010";
    r( 335) := "00111100";
    r( 336) := "01111100";
    r( 337) := "00111100";
    r( 338) := "01111100";
    r( 339) := "00111100";
    r( 340) := "00111110";
    r( 341) := "01000010";
    r( 342) := "01000010";
    r( 343) := "01000010";
    r( 344) := "01000010";
    r( 345) := "00100010";
    r( 346) := "01111110";
    r( 347) := "00111100";
    r( 348) := "00000000";
    r( 349) := "00111100";
    r( 350) := "00001000";
    r( 351) := "00000000";
    r( 352) := "00010000";
    r( 353) := "00000000";
    r( 354) := "01000000";
    r( 355) := "00000000";
    r( 356) := "00000010";
    r( 357) := "00000000";
    r( 358) := "00001100";
    r( 359) := "00000000";
    r( 360) := "01000000";
    r( 361) := "00001000";
    r( 362) := "00000100";
    r( 363) := "01000000";
    r( 364) := "00011000";
    r( 365) := "00000000";
    r( 366) := "00000000";
    r( 367) := "00000000";
    r( 368) := "00000000";
    r( 369) := "00000000";
    r( 370) := "00000000";
    r( 371) := "00000000";
    r( 372) := "00010000";
    r( 373) := "00000000";
    r( 374) := "00000000";
    r( 375) := "00000000";
    r( 376) := "00000000";
    r( 377) := "00000000";
    r( 378) := "00000000";
    r( 379) := "00000100";
    r( 380) := "00001000";
    r( 381) := "00100000";
    r( 382) := "00010100";
    r( 383) := "11111110";
    r( 384) := "00000000";
    r( 385) := "00011000";
    r( 386) := "00011000";
    r( 387) := "00011000";
    r( 388) := "00000000";
    r( 389) := "00000000";
    r( 390) := "00011000";
    r( 391) := "00011000";
    r( 392) := "00011000";
    r( 393) := "00000000";
    r( 394) := "00011000";
    r( 395) := "00000000";
    r( 396) := "00000000";
    r( 397) := "00000000";
    r( 398) := "00000000";
    r( 399) := "00111100";
    r( 400) := "00100100";
    r( 401) := "00000000";
    r( 402) := "00000000";
    r( 403) := "00000000";
    r( 404) := "00000000";
    r( 405) := "00111100";
    r( 406) := "00100100";
    r( 407) := "00000000";
    r( 408) := "00000000";
    r( 409) := "00000000";
    r( 410) := "00000000";
    r( 411) := "00000000";
    r( 412) := "00000000";
    r( 413) := "00000000";
    r( 414) := "00111100";
    r( 415) := "00000000";
    r( 416) := "00000000";
    r( 417) := "00001000";
    r( 418) := "00000000";
    r( 419) := "00001100";
    r( 420) := "00001000";
    r( 421) := "00110000";
    r( 422) := "00001000";
    r( 423) := "00001000";
    r( 424) := "00000100";
    r( 425) := "00010000";
    r( 426) := "00000000";
    r( 427) := "00000000";
    r( 428) := "00000000";
    r( 429) := "00000000";
    r( 430) := "00000000";
    r( 431) := "00000000";
    r( 432) := "00011100";
    r( 433) := "00001000";
    r( 434) := "00011100";
    r( 435) := "00111110";
    r( 436) := "00000100";
    r( 437) := "00111110";
    r( 438) := "00001110";
    r( 439) := "00111110";
    r( 440) := "00011100";
    r( 441) := "00011110";
    r( 442) := "00000000";
    r( 443) := "00000000";
    r( 444) := "00000100";
    r( 445) := "00000000";
    r( 446) := "00100000";
    r( 447) := "00011100";
    r( 448) := "00011100";
    r( 449) := "00001000";
    r( 450) := "00111100";
    r( 451) := "00011100";
    r( 452) := "00111100";
    r( 453) := "00111110";
    r( 454) := "00111110";
    r( 455) := "00011100";
    r( 456) := "00100010";
    r( 457) := "00011100";
    r( 458) := "00000010";
    r( 459) := "00100010";
    r( 460) := "00100000";
    r( 461) := "00100010";
    r( 462) := "00100010";
    r( 463) := "00011100";
    r( 464) := "00111100";
    r( 465) := "00011100";
    r( 466) := "00111100";
    r( 467) := "00011100";
    r( 468) := "00111110";
    r( 469) := "00100010";
    r( 470) := "00100010";
    r( 471) := "00100010";
    r( 472) := "00100010";
    r( 473) := "00100010";
    r( 474) := "00111110";
    r( 475) := "00000000";
    r( 476) := "00010000";
    r( 477) := "00000000";
    r( 478) := "00001000";
    r( 479) := "00000000";
    r( 480) := "00000000";
    r( 481) := "00000000";
    r( 482) := "00100000";
    r( 483) := "00000000";
    r( 484) := "00000010";
    r( 485) := "00000000";
    r( 486) := "00000100";
    r( 487) := "00000000";
    r( 488) := "00100000";
    r( 489) := "00000000";
    r( 490) := "00000000";
    r( 491) := "00100000";
    r( 492) := "00001000";
    r( 493) := "00000000";
    r( 494) := "00000000";
    r( 495) := "00000000";
    r( 496) := "00000000";
    r( 497) := "00000000";
    r( 498) := "00000000";
    r( 499) := "00000000";
    r( 500) := "00000000";
    r( 501) := "00000000";
    r( 502) := "00000000";
    r( 503) := "00000000";
    r( 504) := "00000000";
    r( 505) := "00000000";
    r( 506) := "00000000";
    r( 507) := "00010000";
    r( 508) := "00110110";
    r( 509) := "00110000";
    r( 510) := "00000000";
    r( 511) := "00111110";
    r( 512) := "00000000";
    r( 513) := "00000000";
    r( 514) := "00100100";
    r( 515) := "01000010";
    r( 516) := "10000010";
    r( 517) := "01000010";
    r( 518) := "00001010";
    r( 519) := "00101000";
    r( 520) := "00010000";
    r( 521) := "00001000";
    r( 522) := "00010000";
    r( 523) := "00111000";
    r( 524) := "01010100";
    r( 525) := "00000110";
    r( 526) := "00000010";
    r( 527) := "00000000";
    r( 528) := "11111110";
    r( 529) := "00111000";
    r( 530) := "00111000";
    r( 531) := "00111000";
    r( 532) := "00010000";
    r( 533) := "01000100";
    r( 534) := "01110000";
    r( 535) := "00010000";
    r( 536) := "00100100";
    r( 537) := "00011100";
    r( 538) := "00111000";
    r( 539) := "01111100";
    r( 540) := "01010100";
    r( 541) := "00000100";
    r( 542) := "00010000";
    r( 543) := "00000000";
    r( 544) := "00000000";
    r( 545) := "00001000";
    r( 546) := "00100100";
    r( 547) := "00100100";
    r( 548) := "00011110";
    r( 549) := "01100010";
    r( 550) := "01001000";
    r( 551) := "00001000";
    r( 552) := "00001000";
    r( 553) := "00010000";
    r( 554) := "00101010";
    r( 555) := "00001000";
    r( 556) := "00000000";
    r( 557) := "00000000";
    r( 558) := "00000000";
    r( 559) := "00000010";
    r( 560) := "01000010";
    r( 561) := "00011000";
    r( 562) := "01000010";
    r( 563) := "01000010";
    r( 564) := "00001100";
    r( 565) := "01000000";
    r( 566) := "00100000";
    r( 567) := "01000010";
    r( 568) := "01000010";
    r( 569) := "01000010";
    r( 570) := "00000000";
    r( 571) := "00000000";
    r( 572) := "00001000";
    r( 573) := "00000000";
    r( 574) := "00010000";
    r( 575) := "01000010";
    r( 576) := "00100010";
    r( 577) := "00100100";
    r( 578) := "01000010";
    r( 579) := "01000010";
    r( 580) := "00100010";
    r( 581) := "01000000";
    r( 582) := "01000000";
    r( 583) := "01000010";
    r( 584) := "01000010";
    r( 585) := "00001000";
    r( 586) := "00000100";
    r( 587) := "01000100";
    r( 588) := "01000000";
    r( 589) := "01100110";
    r( 590) := "01100010";
    r( 591) := "01000010";
    r( 592) := "01000010";
    r( 593) := "01000010";
    r( 594) := "01000010";
    r( 595) := "01000010";
    r( 596) := "00001000";
    r( 597) := "01000010";
    r( 598) := "01000010";
    r( 599) := "01000010";
    r( 600) := "01000010";
    r( 601) := "00100010";
    r( 602) := "00000010";
    r( 603) := "00100000";
    r( 604) := "01000000";
    r( 605) := "00000100";
    r( 606) := "00010100";
    r( 607) := "00000000";
    r( 608) := "00001000";
    r( 609) := "00000000";
    r( 610) := "01000000";
    r( 611) := "00000000";
    r( 612) := "00000010";
    r( 613) := "00000000";
    r( 614) := "00010010";
    r( 615) := "00000000";
    r( 616) := "01000000";
    r( 617) := "00000000";
    r( 618) := "00000000";
    r( 619) := "01000000";
    r( 620) := "00001000";
    r( 621) := "00000000";
    r( 622) := "00000000";
    r( 623) := "00000000";
    r( 624) := "00000000";
    r( 625) := "00000000";
    r( 626) := "00000000";
    r( 627) := "00000000";
    r( 628) := "00010000";
    r( 629) := "00000000";
    r( 630) := "00000000";
    r( 631) := "00000000";
    r( 632) := "00000000";
    r( 633) := "00000000";
    r( 634) := "00000000";
    r( 635) := "00001000";
    r( 636) := "00001000";
    r( 637) := "00010000";
    r( 638) := "00101000";
    r( 639) := "11111110";
    r( 640) := "00000000";
    r( 641) := "00011000";
    r( 642) := "00011000";
    r( 643) := "00011000";
    r( 644) := "00000000";
    r( 645) := "00000000";
    r( 646) := "00011000";
    r( 647) := "00011000";
    r( 648) := "00011000";
    r( 649) := "00000000";
    r( 650) := "00011000";
    r( 651) := "00000000";
    r( 652) := "00000000";
    r( 653) := "00000000";
    r( 654) := "00000000";
    r( 655) := "00100100";
    r( 656) := "00100100";
    r( 657) := "00000000";
    r( 658) := "00000000";
    r( 659) := "00000000";
    r( 660) := "00000000";
    r( 661) := "00100100";
    r( 662) := "00100100";
    r( 663) := "00000000";
    r( 664) := "00000000";
    r( 665) := "00000000";
    r( 666) := "00000000";
    r( 667) := "00000000";
    r( 668) := "00000000";
    r( 669) := "00111100";
    r( 670) := "00000000";
    r( 671) := "00000000";
    r( 672) := "00000000";
    r( 673) := "00001000";
    r( 674) := "00010100";
    r( 675) := "00010010";
    r( 676) := "00011110";
    r( 677) := "00110010";
    r( 678) := "00010100";
    r( 679) := "00001000";
    r( 680) := "00001000";
    r( 681) := "00001000";
    r( 682) := "00001000";
    r( 683) := "00001000";
    r( 684) := "00000000";
    r( 685) := "00000000";
    r( 686) := "00000000";
    r( 687) := "00000010";
    r( 688) := "00100010";
    r( 689) := "00011000";
    r( 690) := "00100010";
    r( 691) := "00000010";
    r( 692) := "00001100";
    r( 693) := "00100000";
    r( 694) := "00010000";
    r( 695) := "00000010";
    r( 696) := "00100010";
    r( 697) := "00100010";
    r( 698) := "00000000";
    r( 699) := "00000000";
    r( 700) := "00001000";
    r( 701) := "00000000";
    r( 702) := "00010000";
    r( 703) := "00100010";
    r( 704) := "00100010";
    r( 705) := "00010100";
    r( 706) := "00100010";
    r( 707) := "00100010";
    r( 708) := "00010010";
    r( 709) := "00100000";
    r( 710) := "00100000";
    r( 711) := "00100010";
    r( 712) := "00100010";
    r( 713) := "00001000";
    r( 714) := "00000010";
    r( 715) := "00100100";
    r( 716) := "00100000";
    r( 717) := "00110110";
    r( 718) := "00100010";
    r( 719) := "00100010";
    r( 720) := "00100010";
    r( 721) := "00100010";
    r( 722) := "00100010";
    r( 723) := "00100010";
    r( 724) := "00001000";
    r( 725) := "00100010";
    r( 726) := "00100010";
    r( 727) := "00100010";
    r( 728) := "00100010";
    r( 729) := "00100010";
    r( 730) := "00000010";
    r( 731) := "00001000";
    r( 732) := "00110000";
    r( 733) := "00001000";
    r( 734) := "00011100";
    r( 735) := "00000000";
    r( 736) := "00000000";
    r( 737) := "00000000";
    r( 738) := "00100000";
    r( 739) := "00000000";
    r( 740) := "00000010";
    r( 741) := "00000000";
    r( 742) := "00001000";
    r( 743) := "00000000";
    r( 744) := "00100000";
    r( 745) := "00001000";
    r( 746) := "00001000";
    r( 747) := "00100000";
    r( 748) := "00001000";
    r( 749) := "00000000";
    r( 750) := "00000000";
    r( 751) := "00000000";
    r( 752) := "00000000";
    r( 753) := "00000000";
    r( 754) := "00000000";
    r( 755) := "00000000";
    r( 756) := "00001000";
    r( 757) := "00000000";
    r( 758) := "00000000";
    r( 759) := "00000000";
    r( 760) := "00000000";
    r( 761) := "00000000";
    r( 762) := "00000000";
    r( 763) := "00110000";
    r( 764) := "00110110";
    r( 765) := "00001000";
    r( 766) := "00001000";
    r( 767) := "00111110";
    r( 768) := "00000000";
    r( 769) := "00011000";
    r( 770) := "00100100";
    r( 771) := "01011010";
    r( 772) := "10000010";
    r( 773) := "00100000";
    r( 774) := "00001000";
    r( 775) := "01000100";
    r( 776) := "00100000";
    r( 777) := "00000100";
    r( 778) := "00010000";
    r( 779) := "01010100";
    r( 780) := "00111000";
    r( 781) := "00001110";
    r( 782) := "00000100";
    r( 783) := "00000000";
    r( 784) := "11111110";
    r( 785) := "01111100";
    r( 786) := "01111100";
    r( 787) := "00111000";
    r( 788) := "00010000";
    r( 789) := "00101000";
    r( 790) := "00100000";
    r( 791) := "00000000";
    r( 792) := "00010000";
    r( 793) := "00100000";
    r( 794) := "00010000";
    r( 795) := "00111000";
    r( 796) := "01111100";
    r( 797) := "00011110";
    r( 798) := "00011000";
    r( 799) := "00010000";
    r( 800) := "00000000";
    r( 801) := "00001000";
    r( 802) := "00100100";
    r( 803) := "01111110";
    r( 804) := "00101000";
    r( 805) := "01100100";
    r( 806) := "01001000";
    r( 807) := "00010000";
    r( 808) := "00010000";
    r( 809) := "00001000";
    r( 810) := "00011100";
    r( 811) := "00001000";
    r( 812) := "00000000";
    r( 813) := "00000000";
    r( 814) := "00000000";
    r( 815) := "00000100";
    r( 816) := "01000110";
    r( 817) := "00101000";
    r( 818) := "00000010";
    r( 819) := "00000010";
    r( 820) := "00010100";
    r( 821) := "01111000";
    r( 822) := "01000000";
    r( 823) := "00000100";
    r( 824) := "01000010";
    r( 825) := "01000010";
    r( 826) := "00001000";
    r( 827) := "00001000";
    r( 828) := "00010000";
    r( 829) := "00111100";
    r( 830) := "00001000";
    r( 831) := "00000010";
    r( 832) := "01001010";
    r( 833) := "01000010";
    r( 834) := "01000010";
    r( 835) := "01000000";
    r( 836) := "00100010";
    r( 837) := "01000000";
    r( 838) := "01000000";
    r( 839) := "01000000";
    r( 840) := "01000010";
    r( 841) := "00001000";
    r( 842) := "00000100";
    r( 843) := "01001000";
    r( 844) := "01000000";
    r( 845) := "01011010";
    r( 846) := "01010010";
    r( 847) := "01000010";
    r( 848) := "01000010";
    r( 849) := "01000010";
    r( 850) := "01000010";
    r( 851) := "01000000";
    r( 852) := "00001000";
    r( 853) := "01000010";
    r( 854) := "01000010";
    r( 855) := "01000010";
    r( 856) := "00100100";
    r( 857) := "00100010";
    r( 858) := "00000100";
    r( 859) := "00100000";
    r( 860) := "00100000";
    r( 861) := "00000100";
    r( 862) := "00100010";
    r( 863) := "00000000";
    r( 864) := "00000100";
    r( 865) := "00111000";
    r( 866) := "01011100";
    r( 867) := "00111100";
    r( 868) := "00111010";
    r( 869) := "00111100";
    r( 870) := "00010000";
    r( 871) := "00111010";
    r( 872) := "01011100";
    r( 873) := "00011000";
    r( 874) := "00001100";
    r( 875) := "01000100";
    r( 876) := "00001000";
    r( 877) := "01110100";
    r( 878) := "01111100";
    r( 879) := "00011100";
    r( 880) := "01011100";
    r( 881) := "00111010";
    r( 882) := "01011100";
    r( 883) := "00111110";
    r( 884) := "01111110";
    r( 885) := "01000010";
    r( 886) := "01000010";
    r( 887) := "00100010";
    r( 888) := "01000010";
    r( 889) := "01000010";
    r( 890) := "01111110";
    r( 891) := "00001000";
    r( 892) := "00001000";
    r( 893) := "00010000";
    r( 894) := "00000000";
    r( 895) := "11111110";
    r( 896) := "00000000";
    r( 897) := "00011000";
    r( 898) := "00011000";
    r( 899) := "00011000";
    r( 900) := "00000000";
    r( 901) := "00000000";
    r( 902) := "00011000";
    r( 903) := "00011000";
    r( 904) := "00011000";
    r( 905) := "00000000";
    r( 906) := "00011000";
    r( 907) := "00000000";
    r( 908) := "00000000";
    r( 909) := "00000000";
    r( 910) := "00111100";
    r( 911) := "00100100";
    r( 912) := "00100100";
    r( 913) := "00000000";
    r( 914) := "00000000";
    r( 915) := "00000000";
    r( 916) := "00111100";
    r( 917) := "00100100";
    r( 918) := "00100100";
    r( 919) := "00000000";
    r( 920) := "00000000";
    r( 921) := "00000000";
    r( 922) := "00000000";
    r( 923) := "00000000";
    r( 924) := "00111100";
    r( 925) := "00000000";
    r( 926) := "00000000";
    r( 927) := "00000000";
    r( 928) := "00000000";
    r( 929) := "00001000";
    r( 930) := "00010100";
    r( 931) := "00010000";
    r( 932) := "00101000";
    r( 933) := "00000100";
    r( 934) := "00010100";
    r( 935) := "00010000";
    r( 936) := "00010000";
    r( 937) := "00000100";
    r( 938) := "00101010";
    r( 939) := "00001000";
    r( 940) := "00000000";
    r( 941) := "00000000";
    r( 942) := "00000000";
    r( 943) := "00000100";
    r( 944) := "00110010";
    r( 945) := "00001000";
    r( 946) := "00000010";
    r( 947) := "00000100";
    r( 948) := "00010100";
    r( 949) := "00111100";
    r( 950) := "00100000";
    r( 951) := "00000100";
    r( 952) := "00100010";
    r( 953) := "00100010";
    r( 954) := "00000000";
    r( 955) := "00000000";
    r( 956) := "00010000";
    r( 957) := "00111100";
    r( 958) := "00001000";
    r( 959) := "00000010";
    r( 960) := "00101110";
    r( 961) := "00100010";
    r( 962) := "00100010";
    r( 963) := "00100000";
    r( 964) := "00010010";
    r( 965) := "00100000";
    r( 966) := "00100000";
    r( 967) := "00100000";
    r( 968) := "00100010";
    r( 969) := "00001000";
    r( 970) := "00000010";
    r( 971) := "00101000";
    r( 972) := "00100000";
    r( 973) := "00101010";
    r( 974) := "00110010";
    r( 975) := "00100010";
    r( 976) := "00100010";
    r( 977) := "00100010";
    r( 978) := "00100010";
    r( 979) := "00100000";
    r( 980) := "00001000";
    r( 981) := "00100010";
    r( 982) := "00100010";
    r( 983) := "00100010";
    r( 984) := "00010100";
    r( 985) := "00010100";
    r( 986) := "00000100";
    r( 987) := "00010000";
    r( 988) := "00010000";
    r( 989) := "00000100";
    r( 990) := "00101010";
    r( 991) := "00000000";
    r( 992) := "00000000";
    r( 993) := "00011100";
    r( 994) := "00111100";
    r( 995) := "00011110";
    r( 996) := "00011110";
    r( 997) := "00011100";
    r( 998) := "00001000";
    r( 999) := "00011110";
    r(1000) := "00111100";
    r(1001) := "00000000";
    r(1002) := "00000000";
    r(1003) := "00100100";
    r(1004) := "00001000";
    r(1005) := "00110100";
    r(1006) := "00111100";
    r(1007) := "00011100";
    r(1008) := "00111100";
    r(1009) := "00011110";
    r(1010) := "00101110";
    r(1011) := "00011110";
    r(1012) := "00011100";
    r(1013) := "00100010";
    r(1014) := "00100010";
    r(1015) := "00100010";
    r(1016) := "00100010";
    r(1017) := "00100010";
    r(1018) := "00111110";
    r(1019) := "00010000";
    r(1020) := "00110110";
    r(1021) := "00110000";
    r(1022) := "00000000";
    r(1023) := "00111110";
    r(1024) := "00000000";
    r(1025) := "00100100";
    r(1026) := "00011000";
    r(1027) := "01010010";
    r(1028) := "10010010";
    r(1029) := "00010000";
    r(1030) := "00010000";
    r(1031) := "01000100";
    r(1032) := "01111110";
    r(1033) := "01111110";
    r(1034) := "10010010";
    r(1035) := "10010010";
    r(1036) := "10010010";
    r(1037) := "00011110";
    r(1038) := "00000100";
    r(1039) := "00111110";
    r(1040) := "11111110";
    r(1041) := "11111110";
    r(1042) := "11111110";
    r(1043) := "01010100";
    r(1044) := "01000100";
    r(1045) := "00010000";
    r(1046) := "00100000";
    r(1047) := "01111100";
    r(1048) := "00101000";
    r(1049) := "00100000";
    r(1050) := "00111000";
    r(1051) := "00010000";
    r(1052) := "00111000";
    r(1053) := "00111110";
    r(1054) := "01011100";
    r(1055) := "00111000";
    r(1056) := "00000000";
    r(1057) := "00001000";
    r(1058) := "00000000";
    r(1059) := "00100100";
    r(1060) := "00011100";
    r(1061) := "00001000";
    r(1062) := "00110000";
    r(1063) := "00000000";
    r(1064) := "00010000";
    r(1065) := "00001000";
    r(1066) := "00011100";
    r(1067) := "00111110";
    r(1068) := "00000000";
    r(1069) := "00111100";
    r(1070) := "00000000";
    r(1071) := "00001000";
    r(1072) := "01011010";
    r(1073) := "00001000";
    r(1074) := "00001100";
    r(1075) := "00001100";
    r(1076) := "00100100";
    r(1077) := "00000100";
    r(1078) := "01111100";
    r(1079) := "00001000";
    r(1080) := "00111100";
    r(1081) := "00111110";
    r(1082) := "00000000";
    r(1083) := "00000000";
    r(1084) := "00100000";
    r(1085) := "00000000";
    r(1086) := "00000100";
    r(1087) := "00001100";
    r(1088) := "01010110";
    r(1089) := "01111110";
    r(1090) := "01111100";
    r(1091) := "01000000";
    r(1092) := "00100010";
    r(1093) := "01111000";
    r(1094) := "01111000";
    r(1095) := "01001110";
    r(1096) := "01111110";
    r(1097) := "00001000";
    r(1098) := "00000100";
    r(1099) := "01110000";
    r(1100) := "01000000";
    r(1101) := "01011010";
    r(1102) := "01001010";
    r(1103) := "01000010";
    r(1104) := "01111100";
    r(1105) := "01000010";
    r(1106) := "01111100";
    r(1107) := "00111100";
    r(1108) := "00001000";
    r(1109) := "01000010";
    r(1110) := "00100100";
    r(1111) := "01011010";
    r(1112) := "00011000";
    r(1113) := "00011100";
    r(1114) := "00011000";
    r(1115) := "00100000";
    r(1116) := "00010000";
    r(1117) := "00000100";
    r(1118) := "00000000";
    r(1119) := "00000000";
    r(1120) := "00000000";
    r(1121) := "00000100";
    r(1122) := "01100010";
    r(1123) := "01000000";
    r(1124) := "01000110";
    r(1125) := "01000010";
    r(1126) := "01111100";
    r(1127) := "01000110";
    r(1128) := "01100010";
    r(1129) := "00001000";
    r(1130) := "00000100";
    r(1131) := "01001000";
    r(1132) := "00001000";
    r(1133) := "00101010";
    r(1134) := "00100010";
    r(1135) := "00100010";
    r(1136) := "01100010";
    r(1137) := "01000110";
    r(1138) := "01100010";
    r(1139) := "01000000";
    r(1140) := "00010000";
    r(1141) := "01000010";
    r(1142) := "01000010";
    r(1143) := "00100010";
    r(1144) := "00100100";
    r(1145) := "01000010";
    r(1146) := "00000100";
    r(1147) := "00010000";
    r(1148) := "00001000";
    r(1149) := "00001000";
    r(1150) := "00000000";
    r(1151) := "11111110";
    r(1152) := "11111111";
    r(1153) := "00011000";
    r(1154) := "11111000";
    r(1155) := "00011111";
    r(1156) := "11110000";
    r(1157) := "00001111";
    r(1158) := "11111000";
    r(1159) := "00011111";
    r(1160) := "11111111";
    r(1161) := "11111111";
    r(1162) := "11111111";
    r(1163) := "00000000";
    r(1164) := "00000000";
    r(1165) := "00000000";
    r(1166) := "00100100";
    r(1167) := "00100100";
    r(1168) := "00100100";
    r(1169) := "00000000";
    r(1170) := "00000000";
    r(1171) := "00000000";
    r(1172) := "00100100";
    r(1173) := "00100100";
    r(1174) := "00100100";
    r(1175) := "00000000";
    r(1176) := "00000000";
    r(1177) := "00000000";
    r(1178) := "00000000";
    r(1179) := "00111100";
    r(1180) := "00000000";
    r(1181) := "00000000";
    r(1182) := "00000000";
    r(1183) := "00000000";
    r(1184) := "00000000";
    r(1185) := "00001000";
    r(1186) := "00010100";
    r(1187) := "00011100";
    r(1188) := "00011100";
    r(1189) := "00001000";
    r(1190) := "00011000";
    r(1191) := "00000000";
    r(1192) := "00010000";
    r(1193) := "00000100";
    r(1194) := "00011100";
    r(1195) := "00111110";
    r(1196) := "00000000";
    r(1197) := "00011100";
    r(1198) := "00000000";
    r(1199) := "00001000";
    r(1200) := "00101010";
    r(1201) := "00001000";
    r(1202) := "00001100";
    r(1203) := "00001100";
    r(1204) := "00100100";
    r(1205) := "00000010";
    r(1206) := "00111100";
    r(1207) := "00001000";
    r(1208) := "00011100";
    r(1209) := "00011110";
    r(1210) := "00000000";
    r(1211) := "00001000";
    r(1212) := "00100000";
    r(1213) := "00000000";
    r(1214) := "00000100";
    r(1215) := "00000100";
    r(1216) := "00101010";
    r(1217) := "00100010";
    r(1218) := "00111100";
    r(1219) := "00100000";
    r(1220) := "00010010";
    r(1221) := "00111100";
    r(1222) := "00111100";
    r(1223) := "00100000";
    r(1224) := "00111110";
    r(1225) := "00001000";
    r(1226) := "00000010";
    r(1227) := "00110000";
    r(1228) := "00100000";
    r(1229) := "00101010";
    r(1230) := "00101010";
    r(1231) := "00100010";
    r(1232) := "00111100";
    r(1233) := "00100010";
    r(1234) := "00111100";
    r(1235) := "00011100";
    r(1236) := "00001000";
    r(1237) := "00100010";
    r(1238) := "00010100";
    r(1239) := "00101010";
    r(1240) := "00001000";
    r(1241) := "00001000";
    r(1242) := "00001000";
    r(1243) := "00111110";
    r(1244) := "00010000";
    r(1245) := "00111110";
    r(1246) := "00001000";
    r(1247) := "00000000";
    r(1248) := "00111110";
    r(1249) := "00000010";
    r(1250) := "00100010";
    r(1251) := "00100000";
    r(1252) := "00100010";
    r(1253) := "00100010";
    r(1254) := "00011100";
    r(1255) := "00100010";
    r(1256) := "00100010";
    r(1257) := "00001000";
    r(1258) := "00001000";
    r(1259) := "00101000";
    r(1260) := "00001000";
    r(1261) := "00101010";
    r(1262) := "00100010";
    r(1263) := "00100010";
    r(1264) := "00100010";
    r(1265) := "00100010";
    r(1266) := "00110000";
    r(1267) := "00100000";
    r(1268) := "00001000";
    r(1269) := "00100010";
    r(1270) := "00100010";
    r(1271) := "00100010";
    r(1272) := "00010100";
    r(1273) := "00100010";
    r(1274) := "00000100";
    r(1275) := "00010000";
    r(1276) := "00110110";
    r(1277) := "00001000";
    r(1278) := "00111110";
    r(1279) := "00111110";
    r(1280) := "00001000";
    r(1281) := "01000010";
    r(1282) := "00000000";
    r(1283) := "01011010";
    r(1284) := "10000010";
    r(1285) := "00100000";
    r(1286) := "00010000";
    r(1287) := "01000100";
    r(1288) := "00100000";
    r(1289) := "00000100";
    r(1290) := "01010100";
    r(1291) := "00010000";
    r(1292) := "01010100";
    r(1293) := "00001110";
    r(1294) := "11001000";
    r(1295) := "01010100";
    r(1296) := "01111100";
    r(1297) := "01111100";
    r(1298) := "11111110";
    r(1299) := "11111110";
    r(1300) := "01101100";
    r(1301) := "00101000";
    r(1302) := "00000000";
    r(1303) := "00000000";
    r(1304) := "00010000";
    r(1305) := "00011100";
    r(1306) := "01111100";
    r(1307) := "00111000";
    r(1308) := "00111000";
    r(1309) := "00001100";
    r(1310) := "11011110";
    r(1311) := "00111000";
    r(1312) := "00000000";
    r(1313) := "00000000";
    r(1314) := "00000000";
    r(1315) := "01111110";
    r(1316) := "00001010";
    r(1317) := "00010000";
    r(1318) := "01001010";
    r(1319) := "00000000";
    r(1320) := "00010000";
    r(1321) := "00001000";
    r(1322) := "00011100";
    r(1323) := "00001000";
    r(1324) := "00000000";
    r(1325) := "00000000";
    r(1326) := "00000000";
    r(1327) := "00010000";
    r(1328) := "01100010";
    r(1329) := "00001000";
    r(1330) := "00110000";
    r(1331) := "00000010";
    r(1332) := "01111110";
    r(1333) := "00000010";
    r(1334) := "01000010";
    r(1335) := "00010000";
    r(1336) := "01000010";
    r(1337) := "00000010";
    r(1338) := "00000000";
    r(1339) := "00000000";
    r(1340) := "00010000";
    r(1341) := "00111100";
    r(1342) := "00001000";
    r(1343) := "00010000";
    r(1344) := "01001100";
    r(1345) := "01000010";
    r(1346) := "01000010";
    r(1347) := "01000000";
    r(1348) := "00100010";
    r(1349) := "01000000";
    r(1350) := "01000000";
    r(1351) := "01000010";
    r(1352) := "01000010";
    r(1353) := "00001000";
    r(1354) := "00000100";
    r(1355) := "01001000";
    r(1356) := "01000000";
    r(1357) := "01000010";
    r(1358) := "01000110";
    r(1359) := "01000010";
    r(1360) := "01000000";
    r(1361) := "01001010";
    r(1362) := "01001000";
    r(1363) := "00000010";
    r(1364) := "00001000";
    r(1365) := "01000010";
    r(1366) := "00100100";
    r(1367) := "01011010";
    r(1368) := "00100100";
    r(1369) := "00001000";
    r(1370) := "00100000";
    r(1371) := "00100000";
    r(1372) := "00001000";
    r(1373) := "00000100";
    r(1374) := "00000000";
    r(1375) := "00000000";
    r(1376) := "00000000";
    r(1377) := "00111100";
    r(1378) := "01000010";
    r(1379) := "01000000";
    r(1380) := "01000010";
    r(1381) := "01111110";
    r(1382) := "00010000";
    r(1383) := "01000010";
    r(1384) := "01000010";
    r(1385) := "00001000";
    r(1386) := "00000100";
    r(1387) := "01010000";
    r(1388) := "00001000";
    r(1389) := "00101010";
    r(1390) := "00100010";
    r(1391) := "00100010";
    r(1392) := "01000010";
    r(1393) := "01000010";
    r(1394) := "01000000";
    r(1395) := "00111100";
    r(1396) := "00010000";
    r(1397) := "01000010";
    r(1398) := "01000010";
    r(1399) := "00101010";
    r(1400) := "00011000";
    r(1401) := "01000010";
    r(1402) := "00011000";
    r(1403) := "00001000";
    r(1404) := "00001000";
    r(1405) := "00010000";
    r(1406) := "00000000";
    r(1407) := "11111110";
    r(1408) := "11111111";
    r(1409) := "00011000";
    r(1410) := "11110000";
    r(1411) := "00001111";
    r(1412) := "11111000";
    r(1413) := "00011111";
    r(1414) := "11111000";
    r(1415) := "00011111";
    r(1416) := "11111111";
    r(1417) := "11111111";
    r(1418) := "11111111";
    r(1419) := "00000000";
    r(1420) := "00000000";
    r(1421) := "00111100";
    r(1422) := "00100100";
    r(1423) := "00100100";
    r(1424) := "00100100";
    r(1425) := "00000000";
    r(1426) := "00000000";
    r(1427) := "00111100";
    r(1428) := "00100100";
    r(1429) := "00100100";
    r(1430) := "00100100";
    r(1431) := "00000000";
    r(1432) := "00000000";
    r(1433) := "00000000";
    r(1434) := "00111100";
    r(1435) := "00000000";
    r(1436) := "00000000";
    r(1437) := "00000000";
    r(1438) := "00000000";
    r(1439) := "00000000";
    r(1440) := "00000000";
    r(1441) := "00001000";
    r(1442) := "00000000";
    r(1443) := "00010000";
    r(1444) := "00001010";
    r(1445) := "00010000";
    r(1446) := "00101010";
    r(1447) := "00000000";
    r(1448) := "00010000";
    r(1449) := "00000100";
    r(1450) := "00101010";
    r(1451) := "00001000";
    r(1452) := "00000000";
    r(1453) := "00000000";
    r(1454) := "00000000";
    r(1455) := "00010000";
    r(1456) := "00100110";
    r(1457) := "00001000";
    r(1458) := "00010000";
    r(1459) := "00000010";
    r(1460) := "00111110";
    r(1461) := "00000010";
    r(1462) := "00100010";
    r(1463) := "00010000";
    r(1464) := "00100010";
    r(1465) := "00000010";
    r(1466) := "00010000";
    r(1467) := "00000000";
    r(1468) := "00010000";
    r(1469) := "00111100";
    r(1470) := "00001000";
    r(1471) := "00001000";
    r(1472) := "00101110";
    r(1473) := "00111110";
    r(1474) := "00100010";
    r(1475) := "00100000";
    r(1476) := "00010010";
    r(1477) := "00100000";
    r(1478) := "00100000";
    r(1479) := "00100110";
    r(1480) := "00100010";
    r(1481) := "00001000";
    r(1482) := "00100010";
    r(1483) := "00101000";
    r(1484) := "00100000";
    r(1485) := "00100010";
    r(1486) := "00100110";
    r(1487) := "00100010";
    r(1488) := "00100000";
    r(1489) := "00101010";
    r(1490) := "00101000";
    r(1491) := "00000010";
    r(1492) := "00001000";
    r(1493) := "00100010";
    r(1494) := "00010100";
    r(1495) := "00101010";
    r(1496) := "00010100";
    r(1497) := "00001000";
    r(1498) := "00010000";
    r(1499) := "00010000";
    r(1500) := "00000100";
    r(1501) := "00000100";
    r(1502) := "00001000";
    r(1503) := "00000000";
    r(1504) := "00000000";
    r(1505) := "00011110";
    r(1506) := "00100010";
    r(1507) := "00100000";
    r(1508) := "00100010";
    r(1509) := "00111110";
    r(1510) := "00001000";
    r(1511) := "00100010";
    r(1512) := "00100010";
    r(1513) := "00001000";
    r(1514) := "00001000";
    r(1515) := "00110000";
    r(1516) := "00001000";
    r(1517) := "00101010";
    r(1518) := "00100010";
    r(1519) := "00100010";
    r(1520) := "00100010";
    r(1521) := "00100010";
    r(1522) := "00100000";
    r(1523) := "00011100";
    r(1524) := "00001000";
    r(1525) := "00100010";
    r(1526) := "00010100";
    r(1527) := "00100010";
    r(1528) := "00001000";
    r(1529) := "00100010";
    r(1530) := "00001000";
    r(1531) := "00000010";
    r(1532) := "00110110";
    r(1533) := "00110010";
    r(1534) := "00000000";
    r(1535) := "00111110";
    r(1536) := "00000000";
    r(1537) := "00100100";
    r(1538) := "00000000";
    r(1539) := "01000010";
    r(1540) := "10010010";
    r(1541) := "01000010";
    r(1542) := "00100000";
    r(1543) := "10000010";
    r(1544) := "00010000";
    r(1545) := "00001000";
    r(1546) := "00111000";
    r(1547) := "00010000";
    r(1548) := "00111000";
    r(1549) := "00000110";
    r(1550) := "00101000";
    r(1551) := "00010100";
    r(1552) := "00111000";
    r(1553) := "00111000";
    r(1554) := "01010100";
    r(1555) := "11111110";
    r(1556) := "01010100";
    r(1557) := "01000100";
    r(1558) := "00000000";
    r(1559) := "00010000";
    r(1560) := "01001000";
    r(1561) := "00001000";
    r(1562) := "00111000";
    r(1563) := "00111000";
    r(1564) := "00111000";
    r(1565) := "00011000";
    r(1566) := "01111100";
    r(1567) := "00010000";
    r(1568) := "00000000";
    r(1569) := "00000000";
    r(1570) := "00000000";
    r(1571) := "00100100";
    r(1572) := "00111100";
    r(1573) := "00100110";
    r(1574) := "01000100";
    r(1575) := "00000000";
    r(1576) := "00001000";
    r(1577) := "00010000";
    r(1578) := "00101010";
    r(1579) := "00001000";
    r(1580) := "00000000";
    r(1581) := "00000000";
    r(1582) := "00000000";
    r(1583) := "00100000";
    r(1584) := "01000010";
    r(1585) := "00001000";
    r(1586) := "01000000";
    r(1587) := "01000010";
    r(1588) := "00000100";
    r(1589) := "01000100";
    r(1590) := "01000010";
    r(1591) := "00010000";
    r(1592) := "01000010";
    r(1593) := "00000100";
    r(1594) := "00001000";
    r(1595) := "00001000";
    r(1596) := "00001000";
    r(1597) := "00000000";
    r(1598) := "00010000";
    r(1599) := "00000000";
    r(1600) := "00100000";
    r(1601) := "01000010";
    r(1602) := "01000010";
    r(1603) := "01000010";
    r(1604) := "00100010";
    r(1605) := "01000000";
    r(1606) := "01000000";
    r(1607) := "01000010";
    r(1608) := "01000010";
    r(1609) := "00001000";
    r(1610) := "01000100";
    r(1611) := "01000100";
    r(1612) := "01000000";
    r(1613) := "01000010";
    r(1614) := "01000010";
    r(1615) := "01000010";
    r(1616) := "01000000";
    r(1617) := "01000100";
    r(1618) := "01000100";
    r(1619) := "01000010";
    r(1620) := "00001000";
    r(1621) := "01000010";
    r(1622) := "00011000";
    r(1623) := "01100110";
    r(1624) := "01000010";
    r(1625) := "00001000";
    r(1626) := "01000000";
    r(1627) := "00100000";
    r(1628) := "00000100";
    r(1629) := "00000100";
    r(1630) := "00000000";
    r(1631) := "00000000";
    r(1632) := "00000000";
    r(1633) := "01000100";
    r(1634) := "01100010";
    r(1635) := "01000000";
    r(1636) := "01000110";
    r(1637) := "01000000";
    r(1638) := "00010000";
    r(1639) := "01000110";
    r(1640) := "01000010";
    r(1641) := "00001000";
    r(1642) := "00000100";
    r(1643) := "01101000";
    r(1644) := "00001000";
    r(1645) := "00101010";
    r(1646) := "00100010";
    r(1647) := "00100010";
    r(1648) := "01100010";
    r(1649) := "01000110";
    r(1650) := "01000000";
    r(1651) := "00000010";
    r(1652) := "00010010";
    r(1653) := "01000110";
    r(1654) := "00100100";
    r(1655) := "00101010";
    r(1656) := "00100100";
    r(1657) := "01000110";
    r(1658) := "00100000";
    r(1659) := "00001000";
    r(1660) := "00001000";
    r(1661) := "00010000";
    r(1662) := "00000000";
    r(1663) := "11111110";
    r(1664) := "00000000";
    r(1665) := "00011000";
    r(1666) := "00000000";
    r(1667) := "00000000";
    r(1668) := "00011000";
    r(1669) := "00011000";
    r(1670) := "00011000";
    r(1671) := "00011000";
    r(1672) := "00000000";
    r(1673) := "00011000";
    r(1674) := "00011000";
    r(1675) := "00000000";
    r(1676) := "00000000";
    r(1677) := "00100100";
    r(1678) := "00100100";
    r(1679) := "00100100";
    r(1680) := "00100100";
    r(1681) := "00000000";
    r(1682) := "00000000";
    r(1683) := "00100100";
    r(1684) := "00100100";
    r(1685) := "00100100";
    r(1686) := "00100100";
    r(1687) := "00000000";
    r(1688) := "00000000";
    r(1689) := "00111100";
    r(1690) := "00000000";
    r(1691) := "00000000";
    r(1692) := "00000000";
    r(1693) := "00000000";
    r(1694) := "00000000";
    r(1695) := "00000000";
    r(1696) := "00000000";
    r(1697) := "00000000";
    r(1698) := "00000000";
    r(1699) := "00010000";
    r(1700) := "00111100";
    r(1701) := "00100110";
    r(1702) := "00100100";
    r(1703) := "00000000";
    r(1704) := "00001000";
    r(1705) := "00001000";
    r(1706) := "00001000";
    r(1707) := "00001000";
    r(1708) := "00001000";
    r(1709) := "00000000";
    r(1710) := "00000000";
    r(1711) := "00100000";
    r(1712) := "00100010";
    r(1713) := "00001000";
    r(1714) := "00100000";
    r(1715) := "00100010";
    r(1716) := "00000100";
    r(1717) := "00100010";
    r(1718) := "00100010";
    r(1719) := "00010000";
    r(1720) := "00100010";
    r(1721) := "00000100";
    r(1722) := "00000000";
    r(1723) := "00001000";
    r(1724) := "00001000";
    r(1725) := "00000000";
    r(1726) := "00010000";
    r(1727) := "00000000";
    r(1728) := "00100000";
    r(1729) := "00100010";
    r(1730) := "00100010";
    r(1731) := "00100010";
    r(1732) := "00010010";
    r(1733) := "00100000";
    r(1734) := "00100000";
    r(1735) := "00100010";
    r(1736) := "00100010";
    r(1737) := "00001000";
    r(1738) := "00100010";
    r(1739) := "00100100";
    r(1740) := "00100000";
    r(1741) := "00100010";
    r(1742) := "00100010";
    r(1743) := "00100010";
    r(1744) := "00100000";
    r(1745) := "00100100";
    r(1746) := "00100100";
    r(1747) := "00100010";
    r(1748) := "00001000";
    r(1749) := "00100010";
    r(1750) := "00001000";
    r(1751) := "00101010";
    r(1752) := "00100010";
    r(1753) := "00001000";
    r(1754) := "00100000";
    r(1755) := "00001000";
    r(1756) := "00001010";
    r(1757) := "00001000";
    r(1758) := "00001000";
    r(1759) := "00000000";
    r(1760) := "00000000";
    r(1761) := "00100010";
    r(1762) := "00100010";
    r(1763) := "00100000";
    r(1764) := "00100010";
    r(1765) := "00100000";
    r(1766) := "00001000";
    r(1767) := "00100010";
    r(1768) := "00100010";
    r(1769) := "00001000";
    r(1770) := "00001000";
    r(1771) := "00101000";
    r(1772) := "00001000";
    r(1773) := "00101010";
    r(1774) := "00100010";
    r(1775) := "00100010";
    r(1776) := "00100010";
    r(1777) := "00100010";
    r(1778) := "00100000";
    r(1779) := "00000010";
    r(1780) := "00001000";
    r(1781) := "00100010";
    r(1782) := "00010100";
    r(1783) := "00101010";
    r(1784) := "00010100";
    r(1785) := "00100010";
    r(1786) := "00010000";
    r(1787) := "00000110";
    r(1788) := "00110110";
    r(1789) := "00000110";
    r(1790) := "00001000";
    r(1791) := "00111110";
    r(1792) := "00000000";
    r(1793) := "01100110";
    r(1794) := "00000000";
    r(1795) := "00111100";
    r(1796) := "11111110";
    r(1797) := "11111110";
    r(1798) := "10100000";
    r(1799) := "11111110";
    r(1800) := "00001000";
    r(1801) := "00010000";
    r(1802) := "00010000";
    r(1803) := "00010000";
    r(1804) := "00010000";
    r(1805) := "00000010";
    r(1806) := "00110000";
    r(1807) := "00010100";
    r(1808) := "00010000";
    r(1809) := "00010000";
    r(1810) := "00010000";
    r(1811) := "01010100";
    r(1812) := "01000100";
    r(1813) := "00000000";
    r(1814) := "00000000";
    r(1815) := "00000000";
    r(1816) := "00110000";
    r(1817) := "00000000";
    r(1818) := "01111100";
    r(1819) := "01111100";
    r(1820) := "01111100";
    r(1821) := "00111100";
    r(1822) := "00111000";
    r(1823) := "00111000";
    r(1824) := "00000000";
    r(1825) := "00001000";
    r(1826) := "00000000";
    r(1827) := "00100100";
    r(1828) := "00001000";
    r(1829) := "01000110";
    r(1830) := "00111010";
    r(1831) := "00000000";
    r(1832) := "00000100";
    r(1833) := "00100000";
    r(1834) := "00001000";
    r(1835) := "00000000";
    r(1836) := "00010000";
    r(1837) := "00000000";
    r(1838) := "00010000";
    r(1839) := "01000000";
    r(1840) := "00111100";
    r(1841) := "00111100";
    r(1842) := "01111110";
    r(1843) := "00111100";
    r(1844) := "00000100";
    r(1845) := "00111000";
    r(1846) := "00111100";
    r(1847) := "00010000";
    r(1848) := "00111100";
    r(1849) := "00111000";
    r(1850) := "00000000";
    r(1851) := "00001000";
    r(1852) := "00000100";
    r(1853) := "00000000";
    r(1854) := "00100000";
    r(1855) := "00010000";
    r(1856) := "00011100";
    r(1857) := "01000010";
    r(1858) := "01111100";
    r(1859) := "00111100";
    r(1860) := "01111100";
    r(1861) := "01111110";
    r(1862) := "01000000";
    r(1863) := "00111100";
    r(1864) := "01000010";
    r(1865) := "00011100";
    r(1866) := "00111000";
    r(1867) := "01000010";
    r(1868) := "01111110";
    r(1869) := "01000010";
    r(1870) := "01000010";
    r(1871) := "00111100";
    r(1872) := "01000000";
    r(1873) := "00111010";
    r(1874) := "01000010";
    r(1875) := "00111100";
    r(1876) := "00001000";
    r(1877) := "00111100";
    r(1878) := "00011000";
    r(1879) := "01000010";
    r(1880) := "01000010";
    r(1881) := "00001000";
    r(1882) := "01111110";
    r(1883) := "00111100";
    r(1884) := "00000010";
    r(1885) := "00111100";
    r(1886) := "00000000";
    r(1887) := "00000000";
    r(1888) := "00000000";
    r(1889) := "00111010";
    r(1890) := "01011100";
    r(1891) := "00111100";
    r(1892) := "00111010";
    r(1893) := "00111100";
    r(1894) := "00010000";
    r(1895) := "00111010";
    r(1896) := "01000010";
    r(1897) := "00011100";
    r(1898) := "00000100";
    r(1899) := "01000100";
    r(1900) := "00011100";
    r(1901) := "00101010";
    r(1902) := "00100010";
    r(1903) := "00011100";
    r(1904) := "01011100";
    r(1905) := "00111010";
    r(1906) := "01000000";
    r(1907) := "01111100";
    r(1908) := "00001100";
    r(1909) := "00111010";
    r(1910) := "00011000";
    r(1911) := "00110110";
    r(1912) := "01000010";
    r(1913) := "00111010";
    r(1914) := "01111110";
    r(1915) := "00000100";
    r(1916) := "00001000";
    r(1917) := "00100000";
    r(1918) := "00000000";
    r(1919) := "11111110";
    r(1920) := "00000000";
    r(1921) := "00011000";
    r(1922) := "00000000";
    r(1923) := "00000000";
    r(1924) := "00011000";
    r(1925) := "00011000";
    r(1926) := "00011000";
    r(1927) := "00011000";
    r(1928) := "00000000";
    r(1929) := "00011000";
    r(1930) := "00011000";
    r(1931) := "00000000";
    r(1932) := "00111100";
    r(1933) := "00100100";
    r(1934) := "00100100";
    r(1935) := "00100100";
    r(1936) := "00100100";
    r(1937) := "00000000";
    r(1938) := "00111100";
    r(1939) := "00100100";
    r(1940) := "00100100";
    r(1941) := "00100100";
    r(1942) := "00100100";
    r(1943) := "00000000";
    r(1944) := "00111100";
    r(1945) := "00000000";
    r(1946) := "00000000";
    r(1947) := "00000000";
    r(1948) := "00000000";
    r(1949) := "00000000";
    r(1950) := "00000000";
    r(1951) := "00000000";
    r(1952) := "00000000";
    r(1953) := "00001000";
    r(1954) := "00000000";
    r(1955) := "00101110";
    r(1956) := "00001000";
    r(1957) := "00000110";
    r(1958) := "00011010";
    r(1959) := "00000000";
    r(1960) := "00000100";
    r(1961) := "00010000";
    r(1962) := "00000000";
    r(1963) := "00000000";
    r(1964) := "00001000";
    r(1965) := "00000000";
    r(1966) := "00001000";
    r(1967) := "00000000";
    r(1968) := "00011100";
    r(1969) := "00011100";
    r(1970) := "00111110";
    r(1971) := "00011100";
    r(1972) := "00000100";
    r(1973) := "00011100";
    r(1974) := "00011100";
    r(1975) := "00010000";
    r(1976) := "00011100";
    r(1977) := "00111000";
    r(1978) := "00010000";
    r(1979) := "00001000";
    r(1980) := "00000100";
    r(1981) := "00000000";
    r(1982) := "00100000";
    r(1983) := "00001000";
    r(1984) := "00011100";
    r(1985) := "00100010";
    r(1986) := "00111100";
    r(1987) := "00011100";
    r(1988) := "00111100";
    r(1989) := "00111110";
    r(1990) := "00100000";
    r(1991) := "00011110";
    r(1992) := "00100010";
    r(1993) := "00011100";
    r(1994) := "00011100";
    r(1995) := "00100010";
    r(1996) := "00111110";
    r(1997) := "00100010";
    r(1998) := "00100010";
    r(1999) := "00011100";
    r(2000) := "00100000";
    r(2001) := "00011010";
    r(2002) := "00100010";
    r(2003) := "00011100";
    r(2004) := "00001000";
    r(2005) := "00011100";
    r(2006) := "00001000";
    r(2007) := "00010100";
    r(2008) := "00100010";
    r(2009) := "00001000";
    r(2010) := "00111110";
    r(2011) := "00000000";
    r(2012) := "00000010";
    r(2013) := "00000000";
    r(2014) := "00001000";
    r(2015) := "00111110";
    r(2016) := "00000000";
    r(2017) := "00011110";
    r(2018) := "00111100";
    r(2019) := "00011110";
    r(2020) := "00011110";
    r(2021) := "00011100";
    r(2022) := "00001000";
    r(2023) := "00011110";
    r(2024) := "00100010";
    r(2025) := "00001000";
    r(2026) := "00001000";
    r(2027) := "00100100";
    r(2028) := "00001000";
    r(2029) := "00101010";
    r(2030) := "00100010";
    r(2031) := "00011100";
    r(2032) := "00111100";
    r(2033) := "00011110";
    r(2034) := "00100000";
    r(2035) := "00111100";
    r(2036) := "00000100";
    r(2037) := "00011110";
    r(2038) := "00001000";
    r(2039) := "00010100";
    r(2040) := "00100010";
    r(2041) := "00011110";
    r(2042) := "00111110";
    r(2043) := "00001010";
    r(2044) := "00110110";
    r(2045) := "00001010";
    r(2046) := "00000000";
    r(2047) := "00111110";
    r(2048) := "00000000";
    r(2049) := "00000000";
    r(2050) := "00000000";
    r(2051) := "00000000";
    r(2052) := "00000000";
    r(2053) := "00000000";
    r(2054) := "01000000";
    r(2055) := "00010000";
    r(2056) := "00000000";
    r(2057) := "00000000";
    r(2058) := "00000000";
    r(2059) := "00000000";
    r(2060) := "00000000";
    r(2061) := "00000000";
    r(2062) := "00010000";
    r(2063) := "00000000";
    r(2064) := "00000000";
    r(2065) := "00000000";
    r(2066) := "00000000";
    r(2067) := "00010000";
    r(2068) := "00000000";
    r(2069) := "00000000";
    r(2070) := "00000000";
    r(2071) := "00000000";
    r(2072) := "00000000";
    r(2073) := "00000000";
    r(2074) := "11111110";
    r(2075) := "11111110";
    r(2076) := "11111110";
    r(2077) := "01111110";
    r(2078) := "11111110";
    r(2079) := "01111100";
    r(2080) := "00000000";
    r(2081) := "00000000";
    r(2082) := "00000000";
    r(2083) := "00000000";
    r(2084) := "00000000";
    r(2085) := "00000000";
    r(2086) := "00000000";
    r(2087) := "00000000";
    r(2088) := "00000000";
    r(2089) := "00000000";
    r(2090) := "00000000";
    r(2091) := "00000000";
    r(2092) := "00100000";
    r(2093) := "00000000";
    r(2094) := "00000000";
    r(2095) := "00000000";
    r(2096) := "00000000";
    r(2097) := "00000000";
    r(2098) := "00000000";
    r(2099) := "00000000";
    r(2100) := "00000000";
    r(2101) := "00000000";
    r(2102) := "00000000";
    r(2103) := "00000000";
    r(2104) := "00000000";
    r(2105) := "00000000";
    r(2106) := "00000000";
    r(2107) := "00010000";
    r(2108) := "00000000";
    r(2109) := "00000000";
    r(2110) := "00000000";
    r(2111) := "00000000";
    r(2112) := "00000000";
    r(2113) := "00000000";
    r(2114) := "00000000";
    r(2115) := "00000000";
    r(2116) := "00000000";
    r(2117) := "00000000";
    r(2118) := "00000000";
    r(2119) := "00000000";
    r(2120) := "00000000";
    r(2121) := "00000000";
    r(2122) := "00000000";
    r(2123) := "00000000";
    r(2124) := "00000000";
    r(2125) := "00000000";
    r(2126) := "00000000";
    r(2127) := "00000000";
    r(2128) := "00000000";
    r(2129) := "00000000";
    r(2130) := "00000000";
    r(2131) := "00000000";
    r(2132) := "00000000";
    r(2133) := "00000000";
    r(2134) := "00000000";
    r(2135) := "00000000";
    r(2136) := "00000000";
    r(2137) := "00000000";
    r(2138) := "00000000";
    r(2139) := "00000000";
    r(2140) := "00000000";
    r(2141) := "00000000";
    r(2142) := "00000000";
    r(2143) := "11111111";
    r(2144) := "00000000";
    r(2145) := "00000000";
    r(2146) := "00000000";
    r(2147) := "00000000";
    r(2148) := "00000000";
    r(2149) := "00000000";
    r(2150) := "00000000";
    r(2151) := "00000010";
    r(2152) := "00000000";
    r(2153) := "00000000";
    r(2154) := "01000100";
    r(2155) := "00000000";
    r(2156) := "00000000";
    r(2157) := "00000000";
    r(2158) := "00000000";
    r(2159) := "00000000";
    r(2160) := "01000000";
    r(2161) := "00000010";
    r(2162) := "00000000";
    r(2163) := "00000000";
    r(2164) := "00000000";
    r(2165) := "00000000";
    r(2166) := "00000000";
    r(2167) := "00000000";
    r(2168) := "00000000";
    r(2169) := "00000010";
    r(2170) := "00000000";
    r(2171) := "00000000";
    r(2172) := "00000000";
    r(2173) := "00000000";
    r(2174) := "00000000";
    r(2175) := "11111110";
    r(2176) := "00000000";
    r(2177) := "00011000";
    r(2178) := "00000000";
    r(2179) := "00000000";
    r(2180) := "00011000";
    r(2181) := "00011000";
    r(2182) := "00011000";
    r(2183) := "00011000";
    r(2184) := "00000000";
    r(2185) := "00011000";
    r(2186) := "00011000";
    r(2187) := "00000000";
    r(2188) := "00100100";
    r(2189) := "00100100";
    r(2190) := "00100100";
    r(2191) := "00100100";
    r(2192) := "00100100";
    r(2193) := "00000000";
    r(2194) := "00100100";
    r(2195) := "00100100";
    r(2196) := "00100100";
    r(2197) := "00100100";
    r(2198) := "00100100";
    r(2199) := "00111100";
    r(2200) := "00000000";
    r(2201) := "00000000";
    r(2202) := "00000000";
    r(2203) := "00000000";
    r(2204) := "00000000";
    r(2205) := "00000000";
    r(2206) := "00000000";
    r(2207) := "00000000";
    r(2208) := "00000000";
    r(2209) := "00000000";
    r(2210) := "00000000";
    r(2211) := "00000000";
    r(2212) := "00000000";
    r(2213) := "00000000";
    r(2214) := "00000000";
    r(2215) := "00000000";
    r(2216) := "00000000";
    r(2217) := "00000000";
    r(2218) := "00000000";
    r(2219) := "00000000";
    r(2220) := "00010000";
    r(2221) := "00000000";
    r(2222) := "00000000";
    r(2223) := "00000000";
    r(2224) := "00000000";
    r(2225) := "00000000";
    r(2226) := "00000000";
    r(2227) := "00000000";
    r(2228) := "00000000";
    r(2229) := "00000000";
    r(2230) := "00000000";
    r(2231) := "00000000";
    r(2232) := "00000000";
    r(2233) := "00000000";
    r(2234) := "00000000";
    r(2235) := "00010000";
    r(2236) := "00000000";
    r(2237) := "00000000";
    r(2238) := "00000000";
    r(2239) := "00000000";
    r(2240) := "00000000";
    r(2241) := "00000000";
    r(2242) := "00000000";
    r(2243) := "00000000";
    r(2244) := "00000000";
    r(2245) := "00000000";
    r(2246) := "00000000";
    r(2247) := "00000000";
    r(2248) := "00000000";
    r(2249) := "00000000";
    r(2250) := "00000000";
    r(2251) := "00000000";
    r(2252) := "00000000";
    r(2253) := "00000000";
    r(2254) := "00000000";
    r(2255) := "00000000";
    r(2256) := "00000000";
    r(2257) := "00000000";
    r(2258) := "00000000";
    r(2259) := "00000000";
    r(2260) := "00000000";
    r(2261) := "00000000";
    r(2262) := "00000000";
    r(2263) := "00000000";
    r(2264) := "00000000";
    r(2265) := "00000000";
    r(2266) := "00000000";
    r(2267) := "00000000";
    r(2268) := "00000100";
    r(2269) := "00000000";
    r(2270) := "00000000";
    r(2271) := "00000000";
    r(2272) := "00000000";
    r(2273) := "00000000";
    r(2274) := "00000000";
    r(2275) := "00000000";
    r(2276) := "00000000";
    r(2277) := "00000000";
    r(2278) := "00000000";
    r(2279) := "00000010";
    r(2280) := "00000000";
    r(2281) := "00000000";
    r(2282) := "00001000";
    r(2283) := "00000000";
    r(2284) := "00000000";
    r(2285) := "00000000";
    r(2286) := "00000000";
    r(2287) := "00000000";
    r(2288) := "00100000";
    r(2289) := "00000010";
    r(2290) := "00000000";
    r(2291) := "00000000";
    r(2292) := "00000000";
    r(2293) := "00000000";
    r(2294) := "00000000";
    r(2295) := "00000000";
    r(2296) := "00000000";
    r(2297) := "00000010";
    r(2298) := "00000000";
    r(2299) := "00011110";
    r(2300) := "00000000";
    r(2301) := "00011110";
    r(2302) := "00000000";
    r(2303) := "00000000";
    r(2304) := "00000000";
    r(2305) := "00000000";
    r(2306) := "00000000";
    r(2307) := "00000000";
    r(2308) := "00000000";
    r(2309) := "00000000";
    r(2310) := "00000000";
    r(2311) := "00000000";
    r(2312) := "00000000";
    r(2313) := "00000000";
    r(2314) := "00000000";
    r(2315) := "00000000";
    r(2316) := "00000000";
    r(2317) := "00000000";
    r(2318) := "00000000";
    r(2319) := "00000000";
    r(2320) := "00000000";
    r(2321) := "00000000";
    r(2322) := "00000000";
    r(2323) := "00000000";
    r(2324) := "00000000";
    r(2325) := "00000000";
    r(2326) := "00000000";
    r(2327) := "00000000";
    r(2328) := "00000000";
    r(2329) := "00000000";
    r(2330) := "00000000";
    r(2331) := "00000000";
    r(2332) := "00000000";
    r(2333) := "00000000";
    r(2334) := "00000000";
    r(2335) := "00000000";
    r(2336) := "00000000";
    r(2337) := "00000000";
    r(2338) := "00000000";
    r(2339) := "00000000";
    r(2340) := "00000000";
    r(2341) := "00000000";
    r(2342) := "00000000";
    r(2343) := "00000000";
    r(2344) := "00000000";
    r(2345) := "00000000";
    r(2346) := "00000000";
    r(2347) := "00000000";
    r(2348) := "00000000";
    r(2349) := "00000000";
    r(2350) := "00000000";
    r(2351) := "00000000";
    r(2352) := "00000000";
    r(2353) := "00000000";
    r(2354) := "00000000";
    r(2355) := "00000000";
    r(2356) := "00000000";
    r(2357) := "00000000";
    r(2358) := "00000000";
    r(2359) := "00000000";
    r(2360) := "00000000";
    r(2361) := "00000000";
    r(2362) := "00000000";
    r(2363) := "00000000";
    r(2364) := "00000000";
    r(2365) := "00000000";
    r(2366) := "00000000";
    r(2367) := "00000000";
    r(2368) := "00000000";
    r(2369) := "00000000";
    r(2370) := "00000000";
    r(2371) := "00000000";
    r(2372) := "00000000";
    r(2373) := "00000000";
    r(2374) := "00000000";
    r(2375) := "00000000";
    r(2376) := "00000000";
    r(2377) := "00000000";
    r(2378) := "00000000";
    r(2379) := "00000000";
    r(2380) := "00000000";
    r(2381) := "00000000";
    r(2382) := "00000000";
    r(2383) := "00000000";
    r(2384) := "00000000";
    r(2385) := "00000000";
    r(2386) := "00000000";
    r(2387) := "00000000";
    r(2388) := "00000000";
    r(2389) := "00000000";
    r(2390) := "00000000";
    r(2391) := "00000000";
    r(2392) := "00000000";
    r(2393) := "00000000";
    r(2394) := "00000000";
    r(2395) := "00000000";
    r(2396) := "00000000";
    r(2397) := "00000000";
    r(2398) := "00000000";
    r(2399) := "00000000";
    r(2400) := "00000000";
    r(2401) := "00000000";
    r(2402) := "00000000";
    r(2403) := "00000000";
    r(2404) := "00000000";
    r(2405) := "00000000";
    r(2406) := "00000000";
    r(2407) := "00111100";
    r(2408) := "00000000";
    r(2409) := "00000000";
    r(2410) := "00111000";
    r(2411) := "00000000";
    r(2412) := "00000000";
    r(2413) := "00000000";
    r(2414) := "00000000";
    r(2415) := "00000000";
    r(2416) := "01000000";
    r(2417) := "00000010";
    r(2418) := "00000000";
    r(2419) := "00000000";
    r(2420) := "00000000";
    r(2421) := "00000000";
    r(2422) := "00000000";
    r(2423) := "00000000";
    r(2424) := "00000000";
    r(2425) := "00111100";
    r(2426) := "00000000";
    r(2427) := "00000000";
    r(2428) := "00000000";
    r(2429) := "00000000";
    r(2430) := "00000000";
    r(2431) := "00000000";
    r(2432) := "00000000";
    r(2433) := "00011000";
    r(2434) := "00000000";
    r(2435) := "00000000";
    r(2436) := "00011000";
    r(2437) := "00011000";
    r(2438) := "00011000";
    r(2439) := "00011000";
    r(2440) := "00000000";
    r(2441) := "00011000";
    r(2442) := "00011000";
    r(2443) := "11111111";
    r(2444) := "11111111";
    r(2445) := "11111111";
    r(2446) := "11111111";
    r(2447) := "11111111";
    r(2448) := "11111111";
    r(2449) := "00111100";
    r(2450) := "00100100";
    r(2451) := "00100100";
    r(2452) := "00100100";
    r(2453) := "00100100";
    r(2454) := "00100100";
    r(2455) := "00000000";
    r(2456) := "00000000";
    r(2457) := "00000000";
    r(2458) := "00000000";
    r(2459) := "00000000";
    r(2460) := "00000000";
    r(2461) := "00000000";
    r(2462) := "00000000";
    r(2463) := "00000000";
    r(2464) := "00000000";
    r(2465) := "00000000";
    r(2466) := "00000000";
    r(2467) := "00000000";
    r(2468) := "00000000";
    r(2469) := "00000000";
    r(2470) := "00000000";
    r(2471) := "00000000";
    r(2472) := "00000000";
    r(2473) := "00000000";
    r(2474) := "00000000";
    r(2475) := "00000000";
    r(2476) := "00000000";
    r(2477) := "00000000";
    r(2478) := "00000000";
    r(2479) := "00000000";
    r(2480) := "00000000";
    r(2481) := "00000000";
    r(2482) := "00000000";
    r(2483) := "00000000";
    r(2484) := "00000000";
    r(2485) := "00000000";
    r(2486) := "00000000";
    r(2487) := "00000000";
    r(2488) := "00000000";
    r(2489) := "00000000";
    r(2490) := "00000000";
    r(2491) := "00000000";
    r(2492) := "00000000";
    r(2493) := "00000000";
    r(2494) := "00000000";
    r(2495) := "00000000";
    r(2496) := "00000000";
    r(2497) := "00000000";
    r(2498) := "00000000";
    r(2499) := "00000000";
    r(2500) := "00000000";
    r(2501) := "00000000";
    r(2502) := "00000000";
    r(2503) := "00000000";
    r(2504) := "00000000";
    r(2505) := "00000000";
    r(2506) := "00000000";
    r(2507) := "00000000";
    r(2508) := "00000000";
    r(2509) := "00000000";
    r(2510) := "00000000";
    r(2511) := "00000000";
    r(2512) := "00000000";
    r(2513) := "00000000";
    r(2514) := "00000000";
    r(2515) := "00000000";
    r(2516) := "00000000";
    r(2517) := "00000000";
    r(2518) := "00000000";
    r(2519) := "00000000";
    r(2520) := "00000000";
    r(2521) := "00000000";
    r(2522) := "00000000";
    r(2523) := "00000000";
    r(2524) := "00001010";
    r(2525) := "00000000";
    r(2526) := "00000000";
    r(2527) := "00000000";
    r(2528) := "00000000";
    r(2529) := "00000000";
    r(2530) := "00000000";
    r(2531) := "00000000";
    r(2532) := "00000000";
    r(2533) := "00000000";
    r(2534) := "00000000";
    r(2535) := "00001100";
    r(2536) := "00000000";
    r(2537) := "00000000";
    r(2538) := "00010000";
    r(2539) := "00000000";
    r(2540) := "00000000";
    r(2541) := "00000000";
    r(2542) := "00000000";
    r(2543) := "00000000";
    r(2544) := "00100000";
    r(2545) := "00000010";
    r(2546) := "00000000";
    r(2547) := "00000000";
    r(2548) := "00000000";
    r(2549) := "00000000";
    r(2550) := "00000000";
    r(2551) := "00000000";
    r(2552) := "00000000";
    r(2553) := "00001110";
    r(2554) := "00000000";
    r(2555) := "00000010";
    r(2556) := "00000000";
    r(2557) := "00000010";
    r(2558) := "00000000";
    r(2559) := "00000000";
    return r;
  end init_rom;

  -- Quartus II should notice this and create a .mif file
  signal rom : rom_type := init_rom;

  -- Ensure Quartus II doesn't try to infer an ALTSYNCRAM
  -- as we'd overflow our 26 M4K budget, so instead use LEs
--  attribute ramstyle : string;
--  attribute ramstyle of rom : signal is "logic";

begin

  process ( clk )
  begin
    if rising_edge(clk) then
      q <= rom(to_integer(unsigned(addr)));
    end if;
  end process;

end behavior;
